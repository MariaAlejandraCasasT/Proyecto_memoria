library verilog;
use verilog.vl_types.all;
entity RAM_P_vlg_vec_tst is
end RAM_P_vlg_vec_tst;
