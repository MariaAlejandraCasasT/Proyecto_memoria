library verilog;
use verilog.vl_types.all;
entity PuertosOut_P_vlg_vec_tst is
end PuertosOut_P_vlg_vec_tst;
